/*
Data memory module
Word size: 16 bits, word addressed, size: 1024 bytes. Implemented by reg array in Verilog.
*/
module data_memory()

endmodule
/* 
Branch control unit module
gate-level model required
*/
module branch_control()

endmodule